// inputs are two complex,and each number is 16 bits float

module fft_2_16 (
    input [15:0] i1,i2,
    output [15:0] o1,o2
  );
  
  // this is a temp setting
  parameter W=1

endmodule
